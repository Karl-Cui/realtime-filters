module kernel_lut(kernel, divisor, select);

	output reg [49 * 8 - 1:0] kernel;	// 7x7 8-bit signed coefficients for the chosen kernel in row major order
	output [7:0] divisor;			// 8-bit unsigned normalizing divisor
	input [3:0] select;				// 4-bit kernel selection signal
	
	always @(*) begin
		case (select)
			0: begin  // IDENTITY
					kernel = {	{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00}};
					divisor = 1;
				end
			1: begin  // 3X3 BOX BLUR
					kernel = {	{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h01, 8'h01, 8'h01, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h01, 8'h01, 8'h01, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h01, 8'h01, 8'h01, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00}};
					divisor = 9;
				end
			2: begin  // 5x5 BOX BLUR
					kernel = {{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h00},
								{8'h00, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h00},
								{8'h00, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h00},
								{8'h00, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h00},
								{8'h00, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00}};
					divisor = 25;
				end
			3: begin  // 7x7 BOX BLUR
					kernel = {	{8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01},
								{8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01},
								{8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01},
								{8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01},
								{8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01},
								{8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01},
								{8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01}};
					divisor = 49;
				end
			4: begin  // 3x3 GAUSSIAN BLUR
					kernel = {	{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h01, 8'h02, 8'h01, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h02, 8'h04, 8'h02, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h01, 8'h02, 8'h01, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00}};
					divisor = 16;
				end
			5: begin  // 5x5 GAUSSIAN BLUR
					kernel = {	{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h01, 8'h04, 8'h06, 8'h04, 8'h01, 8'h00},
								{8'h00, 8'h04, 8'h10, 8'h18, 8'h10, 8'h04, 8'h00},
								{8'h00, 8'h06, 8'h18, 8'h23, 8'h18, 8'h06, 8'h00},
								{8'h00, 8'h04, 8'h10, 8'h18, 8'h10, 8'h04, 8'h00},
								{8'h00, 8'h01, 8'h04, 8'h06, 8'h04, 8'h01, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00}};
					divisor = 255;
				end
			6: begin  // 7x7 GAUSSIAN BLUR
					kernel = {	{8'h01, 8'h01, 8'h02, 8'h02, 8'h02, 8'h01, 8'h01},
								{8'h01, 8'h03, 8'h04, 8'h05, 8'h04, 8'h03, 8'h01},
								{8'h02, 8'h04, 8'h07, 8'h08, 8'h07, 8'h04, 8'h02},
								{8'h02, 8'h05, 8'h08, 8'h0A, 8'h08, 8'h05, 8'h02},
								{8'h02, 8'h04, 8'h07, 8'h08, 8'h07, 8'h04, 8'h02},
								{8'h01, 8'h03, 8'h04, 8'h05, 8'h04, 8'h03, 8'h01},
								{8'h01, 8'h01, 8'h02, 8'h02, 8'h02, 8'h01, 8'h01}};
					divisor = 176;
				end
			7: begin  // 3x3 (VERTICAL) SOBEL EDGE DETECTION
					kernel = {	{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'hFF, 8'h00, 8'h01, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'hFE, 8'h00, 8'h02, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'hFF, 8'h00, 8'h01, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00}};
					divisor = 1;
				end
			8: begin  // 3x3 (HORIZONTAL) SOBEL EDGE DETECTION
					kernel = {	{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h01, 8'h02, 8'h01, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'hFF, 8'hFE, 8'hFF, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00}};
					divisor = 1;
				end
			9: begin  // 3x3 SHARPEN
					kernel = {	{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'hFF, 8'h09, 8'hFF, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},
								{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00}};
					divisor = 1;
				end
			default: begin
					kernel = 0;
					divisor = 1;
				end
		endcase
	end
	
endmodule
