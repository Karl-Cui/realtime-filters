module lut(
	 input [1:0] select,
    output reg [44:0] kernel
	 );

    always @(*) begin
      case (select)
        0: kernel = {5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00001, 5'b00000, 5'b00000, 5'b00000, 5'b00000};  // IDENTITY
        1: kernel = {5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001};  // BOX BLUR
        2: kernel = {5'b00001, 5'b00010, 5'b00001, 5'b00010, 5'b00100, 5'b00010, 5'b00001, 5'b00010, 5'b00001};  // GAUSSIAN BLUR
        3: kernel = {5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000};  // SOBEL EDGE DETECTION
//        4: kernel = {5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000};  // SHARPEN
//        5: kernel = {5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000};
//        6: kernel = {5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000};
//        7: kernel = {5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000};
//        default: 
      endcase
    end

endmodule // lut